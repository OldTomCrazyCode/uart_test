//本地测试文件 
module add_test(
    input wire a,
    input wire b,

    output wire c
);
    assign c=a+b;
endmodule

//to push